@00000000
18000000
1820DEAD
A821BEEF
18400000
A8421000
18A00000
A8A50000
E0822800
15000000
D4040800
15000000
9CA50004
15000000
BC050080
15000000
0FFFFFF8
15000000
18A00000
A8A50000
E0822800
15000000
84640000
15000000
9CA50004
15000000
BC050080
15000000
0FFFFFF8
15000000
03FFFFE8
15000000
	 
