@00000000
18000000
18600000
18800000
A8800100
44002000
15000000
	 
