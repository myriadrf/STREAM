@00000000
18000000
1820DEAD
A821BEEF
18400000
A8421000
D4020800
84620000
15000001
15000000
15000000
	 
